--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x: 4
-- 	 network size y: 4
-- 	 Data width: 32
-- 	 Parity: False
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL; 

library work;
use work.type_def_pack.all;

entity network_4x4 is
 generic (DATA_WIDTH: integer := 32; DATA_WIDTH_LV: integer := 11);
port (reset: in  std_logic; 
	clk: in  std_logic; 
	--------------
	RX_L_0: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_0, valid_out_L_0: out std_logic;
	credit_in_L_0, valid_in_L_0: in std_logic;
	TX_L_0: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_1: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_1, valid_out_L_1: out std_logic;
	credit_in_L_1, valid_in_L_1: in std_logic;
	TX_L_1: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_2: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_2, valid_out_L_2: out std_logic;
	credit_in_L_2, valid_in_L_2: in std_logic;
	TX_L_2: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_3: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_3, valid_out_L_3: out std_logic;
	credit_in_L_3, valid_in_L_3: in std_logic;
	TX_L_3: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_4: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_4, valid_out_L_4: out std_logic;
	credit_in_L_4, valid_in_L_4: in std_logic;
	TX_L_4: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_5: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_5, valid_out_L_5: out std_logic;
	credit_in_L_5, valid_in_L_5: in std_logic;
	TX_L_5: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_6: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_6, valid_out_L_6: out std_logic;
	credit_in_L_6, valid_in_L_6: in std_logic;
	TX_L_6: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_7: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_7, valid_out_L_7: out std_logic;
	credit_in_L_7, valid_in_L_7: in std_logic;
	TX_L_7: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_8: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_8, valid_out_L_8: out std_logic;
	credit_in_L_8, valid_in_L_8: in std_logic;
	TX_L_8: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_9: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_9, valid_out_L_9: out std_logic;
	credit_in_L_9, valid_in_L_9: in std_logic;
	TX_L_9: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_10: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_10, valid_out_L_10: out std_logic;
	credit_in_L_10, valid_in_L_10: in std_logic;
	TX_L_10: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_11: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_11, valid_out_L_11: out std_logic;
	credit_in_L_11, valid_in_L_11: in std_logic;
	TX_L_11: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_12: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_12, valid_out_L_12: out std_logic;
	credit_in_L_12, valid_in_L_12: in std_logic;
	TX_L_12: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_13: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_13, valid_out_L_13: out std_logic;
	credit_in_L_13, valid_in_L_13: in std_logic;
	TX_L_13: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_14: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_14, valid_out_L_14: out std_logic;
	credit_in_L_14, valid_in_L_14: in std_logic;
	TX_L_14: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_15: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_15, valid_out_L_15: out std_logic;
	credit_in_L_15, valid_in_L_15: in std_logic;
	TX_L_15: out std_logic_vector (DATA_WIDTH-1 downto 0)

            ); 
end network_4x4; 


architecture behavior of network_4x4 is

--component router_credit_based is
--  generic (
--        DATA_WIDTH: integer := 32; 
--        current_address : integer := 0;
--        Cx_rst : integer := 10;
--        NoC_size: integer := 4
--    );
--    port (
--    reset, clk: in std_logic; 

--    Rxy_reconf: in  std_logic_vector(19 downto 0);
--    Reconfig : in std_logic;
--    RX_N, RX_E, RX_W, RX_S, RX_L : in std_logic_vector (DATA_WIDTH-1 downto 0); 
--    credit_in_N, credit_in_E, credit_in_W, credit_in_S, credit_in_L: in std_logic;
--    valid_in_N, valid_in_E, valid_in_W, valid_in_S, valid_in_L : in std_logic;

--    valid_out_N, valid_out_E, valid_out_W, valid_out_S, valid_out_L : out std_logic;
--    credit_out_N, credit_out_E, credit_out_W, credit_out_S, credit_out_L: out std_logic;

--    TX_N, TX_E, TX_W, TX_S, TX_L: out std_logic_vector (DATA_WIDTH-1 downto 0)
--    ); 
--end component; 

component router_credit_based is
	generic (
        DATA_WIDTH: integer := 32;
        current_address : integer := 0;
        NoC_size: integer := 4; 

        routing_table_bits_local: t_tata := (
            0 =>    "0000",
            1 =>    "0000",
            2 =>    "0000",
            3 =>    "0000",
            4 =>    "0000",
            5 =>    "0000",
            6 =>    "0000",
            7 =>    "0000",
            8 =>    "0000",
            9 =>    "0000",
            10 =>   "0000",
            11 =>   "0000",
            12 =>   "0000",
            13 =>   "0000",
            14 =>   "0000",
            15 =>   "0100"
        ); 

        routing_table_bits_north: t_tata := (
            0 =>    "0000",
            1 =>    "0000",
            2 =>    "0000",
            3 =>    "0000",
            4 =>    "0000",
            5 =>    "0000",
            6 =>    "0000",
            7 =>    "0000",
            8 =>    "0000",
            9 =>    "0000",
            10 =>   "0000",
            11 =>   "0000",
            12 =>   "0000",
            13 =>   "0000",
            14 =>   "0000",
            15 =>   "0100"
        ); 

        routing_table_bits_east: t_tata := (
            0 =>    "0000",
            1 =>    "0000",
            2 =>    "0000",
            3 =>    "0000",
            4 =>    "0000",
            5 =>    "0000",
            6 =>    "0000",
            7 =>    "0000",
            8 =>    "0000",
            9 =>    "0000",
            10 =>   "0000",
            11 =>   "0000",
            12 =>   "0000",
            13 =>   "0000",
            14 =>   "0000",
            15 =>   "0100"
        ); 

        routing_table_bits_west: t_tata := (
            0 =>    "0000",
            1 =>    "0000",
            2 =>    "0000",
            3 =>    "0000",
            4 =>    "0000",
            5 =>    "0000",
            6 =>    "0000",
            7 =>    "0000",
            8 =>    "0000",
            9 =>    "0000",
            10 =>   "0000",
            11 =>   "0000",
            12 =>   "0000",
            13 =>   "0000",
            14 =>   "0000",
            15 =>   "0100"
        );

        routing_table_bits_south: t_tata := (
            0 =>    "0000",
            1 =>    "0000",
            2 =>    "0000",
            3 =>    "0000",
            4 =>    "0000",
            5 =>    "0000",
            6 =>    "0000",
            7 =>    "0000",
            8 =>    "0000",
            9 =>    "0000",
            10 =>   "0000",
            11 =>   "0000",
            12 =>   "0000",
            13 =>   "0000",
            14 =>   "0000",
            15 =>   "0100"
        )
    );
    port (
    reset, clk: in std_logic;

    RX_N, RX_E, RX_W, RX_S, RX_L : in std_logic_vector (DATA_WIDTH-1 downto 0);

    credit_in_N, credit_in_E, credit_in_W, credit_in_S, credit_in_L: in std_logic;
    valid_in_N, valid_in_E, valid_in_W, valid_in_S, valid_in_L : in std_logic;

    valid_out_N, valid_out_E, valid_out_W, valid_out_S, valid_out_L : out std_logic;
    credit_out_N, credit_out_E, credit_out_W, credit_out_S, credit_out_L: out std_logic;

    TX_N, TX_E, TX_W, TX_S, TX_L: out std_logic_vector (DATA_WIDTH-1 downto 0)
    );
end component;



-- generating bulk signals. not all of them are used in the design...
	signal credit_out_N_0, credit_out_E_0, credit_out_W_0, credit_out_S_0: std_logic;
	signal credit_out_N_1, credit_out_E_1, credit_out_W_1, credit_out_S_1: std_logic;
	signal credit_out_N_2, credit_out_E_2, credit_out_W_2, credit_out_S_2: std_logic;
	signal credit_out_N_3, credit_out_E_3, credit_out_W_3, credit_out_S_3: std_logic;
	signal credit_out_N_4, credit_out_E_4, credit_out_W_4, credit_out_S_4: std_logic;
	signal credit_out_N_5, credit_out_E_5, credit_out_W_5, credit_out_S_5: std_logic;
	signal credit_out_N_6, credit_out_E_6, credit_out_W_6, credit_out_S_6: std_logic;
	signal credit_out_N_7, credit_out_E_7, credit_out_W_7, credit_out_S_7: std_logic;
	signal credit_out_N_8, credit_out_E_8, credit_out_W_8, credit_out_S_8: std_logic;
	signal credit_out_N_9, credit_out_E_9, credit_out_W_9, credit_out_S_9: std_logic;
	signal credit_out_N_10, credit_out_E_10, credit_out_W_10, credit_out_S_10: std_logic;
	signal credit_out_N_11, credit_out_E_11, credit_out_W_11, credit_out_S_11: std_logic;
	signal credit_out_N_12, credit_out_E_12, credit_out_W_12, credit_out_S_12: std_logic;
	signal credit_out_N_13, credit_out_E_13, credit_out_W_13, credit_out_S_13: std_logic;
	signal credit_out_N_14, credit_out_E_14, credit_out_W_14, credit_out_S_14: std_logic;
	signal credit_out_N_15, credit_out_E_15, credit_out_W_15, credit_out_S_15: std_logic;

	signal credit_in_N_0, credit_in_E_0, credit_in_W_0, credit_in_S_0: std_logic;
	signal credit_in_N_1, credit_in_E_1, credit_in_W_1, credit_in_S_1: std_logic;
	signal credit_in_N_2, credit_in_E_2, credit_in_W_2, credit_in_S_2: std_logic;
	signal credit_in_N_3, credit_in_E_3, credit_in_W_3, credit_in_S_3: std_logic;
	signal credit_in_N_4, credit_in_E_4, credit_in_W_4, credit_in_S_4: std_logic;
	signal credit_in_N_5, credit_in_E_5, credit_in_W_5, credit_in_S_5: std_logic;
	signal credit_in_N_6, credit_in_E_6, credit_in_W_6, credit_in_S_6: std_logic;
	signal credit_in_N_7, credit_in_E_7, credit_in_W_7, credit_in_S_7: std_logic;
	signal credit_in_N_8, credit_in_E_8, credit_in_W_8, credit_in_S_8: std_logic;
	signal credit_in_N_9, credit_in_E_9, credit_in_W_9, credit_in_S_9: std_logic;
	signal credit_in_N_10, credit_in_E_10, credit_in_W_10, credit_in_S_10: std_logic;
	signal credit_in_N_11, credit_in_E_11, credit_in_W_11, credit_in_S_11: std_logic;
	signal credit_in_N_12, credit_in_E_12, credit_in_W_12, credit_in_S_12: std_logic;
	signal credit_in_N_13, credit_in_E_13, credit_in_W_13, credit_in_S_13: std_logic;
	signal credit_in_N_14, credit_in_E_14, credit_in_W_14, credit_in_S_14: std_logic;
	signal credit_in_N_15, credit_in_E_15, credit_in_W_15, credit_in_S_15: std_logic;

	signal RX_N_0, RX_E_0, RX_W_0, RX_S_0 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_1, RX_E_1, RX_W_1, RX_S_1 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_2, RX_E_2, RX_W_2, RX_S_2 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_3, RX_E_3, RX_W_3, RX_S_3 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_4, RX_E_4, RX_W_4, RX_S_4 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_5, RX_E_5, RX_W_5, RX_S_5 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_6, RX_E_6, RX_W_6, RX_S_6 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_7, RX_E_7, RX_W_7, RX_S_7 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_8, RX_E_8, RX_W_8, RX_S_8 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_9, RX_E_9, RX_W_9, RX_S_9 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_10, RX_E_10, RX_W_10, RX_S_10 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_11, RX_E_11, RX_W_11, RX_S_11 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_12, RX_E_12, RX_W_12, RX_S_12 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_13, RX_E_13, RX_W_13, RX_S_13 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_14, RX_E_14, RX_W_14, RX_S_14 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_15, RX_E_15, RX_W_15, RX_S_15 : std_logic_vector (DATA_WIDTH-1 downto 0);

	signal valid_out_N_0, valid_out_E_0, valid_out_W_0, valid_out_S_0: std_logic;
	signal valid_out_N_1, valid_out_E_1, valid_out_W_1, valid_out_S_1: std_logic;
	signal valid_out_N_2, valid_out_E_2, valid_out_W_2, valid_out_S_2: std_logic;
	signal valid_out_N_3, valid_out_E_3, valid_out_W_3, valid_out_S_3: std_logic;
	signal valid_out_N_4, valid_out_E_4, valid_out_W_4, valid_out_S_4: std_logic;
	signal valid_out_N_5, valid_out_E_5, valid_out_W_5, valid_out_S_5: std_logic;
	signal valid_out_N_6, valid_out_E_6, valid_out_W_6, valid_out_S_6: std_logic;
	signal valid_out_N_7, valid_out_E_7, valid_out_W_7, valid_out_S_7: std_logic;
	signal valid_out_N_8, valid_out_E_8, valid_out_W_8, valid_out_S_8: std_logic;
	signal valid_out_N_9, valid_out_E_9, valid_out_W_9, valid_out_S_9: std_logic;
	signal valid_out_N_10, valid_out_E_10, valid_out_W_10, valid_out_S_10: std_logic;
	signal valid_out_N_11, valid_out_E_11, valid_out_W_11, valid_out_S_11: std_logic;
	signal valid_out_N_12, valid_out_E_12, valid_out_W_12, valid_out_S_12: std_logic;
	signal valid_out_N_13, valid_out_E_13, valid_out_W_13, valid_out_S_13: std_logic;
	signal valid_out_N_14, valid_out_E_14, valid_out_W_14, valid_out_S_14: std_logic;
	signal valid_out_N_15, valid_out_E_15, valid_out_W_15, valid_out_S_15: std_logic;

	signal valid_in_N_0, valid_in_E_0, valid_in_W_0, valid_in_S_0: std_logic;
	signal valid_in_N_1, valid_in_E_1, valid_in_W_1, valid_in_S_1: std_logic;
	signal valid_in_N_2, valid_in_E_2, valid_in_W_2, valid_in_S_2: std_logic;
	signal valid_in_N_3, valid_in_E_3, valid_in_W_3, valid_in_S_3: std_logic;
	signal valid_in_N_4, valid_in_E_4, valid_in_W_4, valid_in_S_4: std_logic;
	signal valid_in_N_5, valid_in_E_5, valid_in_W_5, valid_in_S_5: std_logic;
	signal valid_in_N_6, valid_in_E_6, valid_in_W_6, valid_in_S_6: std_logic;
	signal valid_in_N_7, valid_in_E_7, valid_in_W_7, valid_in_S_7: std_logic;
	signal valid_in_N_8, valid_in_E_8, valid_in_W_8, valid_in_S_8: std_logic;
	signal valid_in_N_9, valid_in_E_9, valid_in_W_9, valid_in_S_9: std_logic;
	signal valid_in_N_10, valid_in_E_10, valid_in_W_10, valid_in_S_10: std_logic;
	signal valid_in_N_11, valid_in_E_11, valid_in_W_11, valid_in_S_11: std_logic;
	signal valid_in_N_12, valid_in_E_12, valid_in_W_12, valid_in_S_12: std_logic;
	signal valid_in_N_13, valid_in_E_13, valid_in_W_13, valid_in_S_13: std_logic;
	signal valid_in_N_14, valid_in_E_14, valid_in_W_14, valid_in_S_14: std_logic;
	signal valid_in_N_15, valid_in_E_15, valid_in_W_15, valid_in_S_15: std_logic;

	signal TX_N_0, TX_E_0, TX_W_0, TX_S_0 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_1, TX_E_1, TX_W_1, TX_S_1 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_2, TX_E_2, TX_W_2, TX_S_2 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_3, TX_E_3, TX_W_3, TX_S_3 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_4, TX_E_4, TX_W_4, TX_S_4 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_5, TX_E_5, TX_W_5, TX_S_5 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_6, TX_E_6, TX_W_6, TX_S_6 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_7, TX_E_7, TX_W_7, TX_S_7 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_8, TX_E_8, TX_W_8, TX_S_8 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_9, TX_E_9, TX_W_9, TX_S_9 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_10, TX_E_10, TX_W_10, TX_S_10 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_11, TX_E_11, TX_W_11, TX_S_11 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_12, TX_E_12, TX_W_12, TX_S_12 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_13, TX_E_13, TX_W_13, TX_S_13 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_14, TX_E_14, TX_W_14, TX_S_14 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_15, TX_E_15, TX_W_15, TX_S_15 : std_logic_vector (DATA_WIDTH-1 downto 0);

-- Node 0
constant routing_table_bits_0: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0000",
		2 => "0000",
		3 => "0000",
		4 => "0000",
		5 => "0000",
		6 => "0000",
		7 => "0000",
		8 => "0000",
		9 => "0000",
		10 => "0000",
		11 => "0000",
		12 => "0000",
		13 => "0000",
		14 => "0000",
		15 => "0100",
	-- north
		16 => "0000",
		17 => "0000",
		18 => "0000",
		19 => "0000",
		20 => "0000",
		21 => "0000",
		22 => "0000",
		23 => "0000",
		24 => "0000",
		25 => "0000",
		26 => "0000",
		27 => "0000",
		28 => "0000",
		29 => "0000",
		30 => "0000",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "0000",
		34 => "0000",
		35 => "0000",
		36 => "0000",
		37 => "0000",
		38 => "0000",
		39 => "0000",
		40 => "0000",
		41 => "0000",
		42 => "0000",
		43 => "0000",
		44 => "0000",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 1
constant routing_table_bits_1: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0000",
		2 => "0001",
		3 => "0000",
		4 => "0001",
		5 => "0001",
		6 => "0001",
		7 => "0001",
		8 => "0001",
		9 => "0001",
		10 => "0001",
		11 => "0001",
		12 => "0001",
		13 => "0001",
		14 => "0001",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0000",
		18 => "0000",
		19 => "0000",
		20 => "0000",
		21 => "0000",
		22 => "0000",
		23 => "0000",
		24 => "0000",
		25 => "0000",
		26 => "0000",
		27 => "0000",
		28 => "0000",
		29 => "0000",
		30 => "0000",
		31 => "0000",
	-- east
		32 => "0010",
		33 => "0000",
		34 => "0000",
		35 => "0000",
		36 => "0000",
		37 => "0000",
		38 => "0000",
		39 => "0000",
		40 => "0000",
		41 => "0000",
		42 => "0000",
		43 => "0000",
		44 => "0000",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0100",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 2
constant routing_table_bits_2: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0001",
		2 => "0000",
		3 => "0000",
		4 => "0001",
		5 => "0001",
		6 => "0001",
		7 => "0001",
		8 => "0001",
		9 => "0001",
		10 => "0001",
		11 => "0001",
		12 => "0001",
		13 => "0001",
		14 => "0001",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0000",
		18 => "0000",
		19 => "0000",
		20 => "0000",
		21 => "0000",
		22 => "0000",
		23 => "0000",
		24 => "0000",
		25 => "0000",
		26 => "0000",
		27 => "0000",
		28 => "0000",
		29 => "0000",
		30 => "0000",
		31 => "0000",
	-- east
		32 => "0010",
		33 => "0000",
		34 => "0000",
		35 => "0000",
		36 => "0000",
		37 => "0000",
		38 => "0000",
		39 => "0000",
		40 => "0000",
		41 => "0000",
		42 => "0000",
		43 => "0000",
		44 => "0000",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0100",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 3
constant routing_table_bits_3: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0000",
		2 => "0000",
		3 => "0000",
		4 => "0000",
		5 => "0000",
		6 => "0000",
		7 => "0000",
		8 => "0000",
		9 => "0000",
		10 => "0000",
		11 => "0000",
		12 => "0000",
		13 => "0000",
		14 => "0000",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0000",
		18 => "0000",
		19 => "0000",
		20 => "0000",
		21 => "0000",
		22 => "0000",
		23 => "0000",
		24 => "0000",
		25 => "0000",
		26 => "0000",
		27 => "0000",
		28 => "0000",
		29 => "0000",
		30 => "0000",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "0000",
		34 => "0000",
		35 => "0000",
		36 => "0000",
		37 => "0000",
		38 => "0000",
		39 => "0000",
		40 => "0000",
		41 => "0000",
		42 => "0000",
		43 => "0000",
		44 => "0000",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0001",
	-- south
		64 => "0010",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 4
constant routing_table_bits_4: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0101",
		2 => "0101",
		3 => "0000",
		4 => "0000",
		5 => "0101",
		6 => "0101",
		7 => "0100",
		8 => "0101",
		9 => "0101",
		10 => "0101",
		11 => "0101",
		12 => "0101",
		13 => "0101",
		14 => "0101",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0000",
		18 => "0000",
		19 => "0000",
		20 => "0000",
		21 => "0000",
		22 => "0000",
		23 => "0000",
		24 => "0000",
		25 => "0000",
		26 => "0000",
		27 => "0000",
		28 => "0000",
		29 => "0000",
		30 => "0000",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "0001",
		34 => "0001",
		35 => "0000",
		36 => "0000",
		37 => "0001",
		38 => "0001",
		39 => "0000",
		40 => "0001",
		41 => "0001",
		42 => "0001",
		43 => "0001",
		44 => "0001",
		45 => "0001",
		46 => "0001",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 5
constant routing_table_bits_5: t_tata_long := (
	-- local
		0 => "0000",
		1 => "1110",
		2 => "0111",
		3 => "0000",
		4 => "0111",
		5 => "0000",
		6 => "0111",
		7 => "0100",
		8 => "0111",
		9 => "0111",
		10 => "0111",
		11 => "0111",
		12 => "0111",
		13 => "0111",
		14 => "0111",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0111",
		18 => "0111",
		19 => "0000",
		20 => "0111",
		21 => "0000",
		22 => "0111",
		23 => "0100",
		24 => "0111",
		25 => "0111",
		26 => "0111",
		27 => "0111",
		28 => "0111",
		29 => "0111",
		30 => "0111",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "1010",
		34 => "0011",
		35 => "0000",
		36 => "0011",
		37 => "0000",
		38 => "0011",
		39 => "0000",
		40 => "0011",
		41 => "0011",
		42 => "0011",
		43 => "0011",
		44 => "0011",
		45 => "0011",
		46 => "0011",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "1100",
		50 => "0101",
		51 => "0000",
		52 => "0101",
		53 => "0000",
		54 => "0101",
		55 => "0100",
		56 => "0101",
		57 => "0101",
		58 => "0101",
		59 => "0101",
		60 => "0101",
		61 => "0101",
		62 => "0101",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "1000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 6
constant routing_table_bits_6: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0011",
		2 => "0011",
		3 => "0000",
		4 => "0011",
		5 => "0011",
		6 => "0000",
		7 => "0100",
		8 => "0011",
		9 => "0011",
		10 => "0011",
		11 => "0011",
		12 => "0011",
		13 => "0011",
		14 => "0011",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0011",
		18 => "0011",
		19 => "0000",
		20 => "0011",
		21 => "0011",
		22 => "0000",
		23 => "0100",
		24 => "0011",
		25 => "0011",
		26 => "0011",
		27 => "0011",
		28 => "0011",
		29 => "0011",
		30 => "0011",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "0011",
		34 => "0011",
		35 => "0000",
		36 => "0011",
		37 => "0011",
		38 => "0000",
		39 => "0000",
		40 => "0011",
		41 => "0011",
		42 => "0011",
		43 => "0011",
		44 => "0011",
		45 => "0011",
		46 => "0011",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0001",
		50 => "0001",
		51 => "0000",
		52 => "0001",
		53 => "0001",
		54 => "0000",
		55 => "0100",
		56 => "0001",
		57 => "0001",
		58 => "0001",
		59 => "0001",
		60 => "0001",
		61 => "0001",
		62 => "0001",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "1000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 7
constant routing_table_bits_7: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0010",
		2 => "0010",
		3 => "0000",
		4 => "0010",
		5 => "0010",
		6 => "0010",
		7 => "0000",
		8 => "0010",
		9 => "0010",
		10 => "0010",
		11 => "0010",
		12 => "0010",
		13 => "0010",
		14 => "0010",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0000",
		18 => "0000",
		19 => "0000",
		20 => "0000",
		21 => "0000",
		22 => "0000",
		23 => "0000",
		24 => "0000",
		25 => "0000",
		26 => "0000",
		27 => "0000",
		28 => "0000",
		29 => "0000",
		30 => "0000",
		31 => "0001",
	-- east
		32 => "0000",
		33 => "0000",
		34 => "0000",
		35 => "0000",
		36 => "0000",
		37 => "0000",
		38 => "0000",
		39 => "0000",
		40 => "0000",
		41 => "0000",
		42 => "0000",
		43 => "0000",
		44 => "0000",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0000",
	-- south
		64 => "1000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 8
constant routing_table_bits_8: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0101",
		2 => "0101",
		3 => "0000",
		4 => "1100",
		5 => "0101",
		6 => "0101",
		7 => "0000",
		8 => "0000",
		9 => "0101",
		10 => "0101",
		11 => "0100",
		12 => "0101",
		13 => "0101",
		14 => "0101",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0101",
		18 => "0101",
		19 => "0000",
		20 => "0100",
		21 => "0101",
		22 => "0101",
		23 => "0000",
		24 => "0000",
		25 => "0101",
		26 => "0101",
		27 => "0100",
		28 => "0101",
		29 => "0101",
		30 => "0101",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "0001",
		34 => "0001",
		35 => "0000",
		36 => "1000",
		37 => "0001",
		38 => "0001",
		39 => "0000",
		40 => "0000",
		41 => "0001",
		42 => "0001",
		43 => "0000",
		44 => "0001",
		45 => "0001",
		46 => "0001",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "1000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 9
constant routing_table_bits_9: t_tata_long := (
	-- local
		0 => "0000",
		1 => "1110",
		2 => "0111",
		3 => "0000",
		4 => "0111",
		5 => "1110",
		6 => "0111",
		7 => "0000",
		8 => "0111",
		9 => "0000",
		10 => "0111",
		11 => "0100",
		12 => "0111",
		13 => "0111",
		14 => "0111",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0110",
		18 => "0111",
		19 => "0000",
		20 => "0111",
		21 => "0110",
		22 => "0111",
		23 => "0000",
		24 => "0111",
		25 => "0000",
		26 => "0111",
		27 => "0100",
		28 => "0111",
		29 => "0111",
		30 => "0111",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "1010",
		34 => "0011",
		35 => "0000",
		36 => "0011",
		37 => "1010",
		38 => "0011",
		39 => "0000",
		40 => "0011",
		41 => "0000",
		42 => "0011",
		43 => "0000",
		44 => "0011",
		45 => "0011",
		46 => "0011",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "1100",
		50 => "0101",
		51 => "0000",
		52 => "0101",
		53 => "1100",
		54 => "0101",
		55 => "0000",
		56 => "0101",
		57 => "0000",
		58 => "0101",
		59 => "0100",
		60 => "0101",
		61 => "0101",
		62 => "0101",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "1000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "1000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 10
constant routing_table_bits_10: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0011",
		2 => "1010",
		3 => "0000",
		4 => "0011",
		5 => "0011",
		6 => "1010",
		7 => "0000",
		8 => "0011",
		9 => "0011",
		10 => "0000",
		11 => "0100",
		12 => "0011",
		13 => "0011",
		14 => "0011",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0011",
		18 => "0010",
		19 => "0000",
		20 => "0011",
		21 => "0011",
		22 => "0010",
		23 => "0000",
		24 => "0011",
		25 => "0011",
		26 => "0000",
		27 => "0100",
		28 => "0011",
		29 => "0011",
		30 => "0011",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "0011",
		34 => "1010",
		35 => "0000",
		36 => "0011",
		37 => "0011",
		38 => "1010",
		39 => "0000",
		40 => "0011",
		41 => "0011",
		42 => "0000",
		43 => "0000",
		44 => "0011",
		45 => "0011",
		46 => "0011",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0001",
		50 => "1000",
		51 => "0000",
		52 => "0001",
		53 => "0001",
		54 => "1000",
		55 => "0000",
		56 => "0001",
		57 => "0001",
		58 => "0000",
		59 => "0100",
		60 => "0001",
		61 => "0001",
		62 => "0001",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "1000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "1000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 11
constant routing_table_bits_11: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0010",
		2 => "0010",
		3 => "0000",
		4 => "0010",
		5 => "0010",
		6 => "0010",
		7 => "0000",
		8 => "0010",
		9 => "0010",
		10 => "0010",
		11 => "0000",
		12 => "0010",
		13 => "0010",
		14 => "0010",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0000",
		18 => "0000",
		19 => "0000",
		20 => "0000",
		21 => "0000",
		22 => "0000",
		23 => "0000",
		24 => "0000",
		25 => "0000",
		26 => "0000",
		27 => "0000",
		28 => "0000",
		29 => "0000",
		30 => "0000",
		31 => "0001",
	-- east
		32 => "0000",
		33 => "0000",
		34 => "0000",
		35 => "0000",
		36 => "0000",
		37 => "0000",
		38 => "0000",
		39 => "0000",
		40 => "0000",
		41 => "0000",
		42 => "0000",
		43 => "0000",
		44 => "0000",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0000",
	-- south
		64 => "1000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 12
constant routing_table_bits_12: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0100",
		2 => "0100",
		3 => "0000",
		4 => "1000",
		5 => "0100",
		6 => "0100",
		7 => "0000",
		8 => "1000",
		9 => "0100",
		10 => "0100",
		11 => "0000",
		12 => "0000",
		13 => "0100",
		14 => "0100",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0100",
		18 => "0100",
		19 => "0000",
		20 => "0000",
		21 => "0100",
		22 => "0100",
		23 => "0000",
		24 => "0000",
		25 => "0100",
		26 => "0100",
		27 => "0000",
		28 => "0000",
		29 => "0100",
		30 => "0100",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "0000",
		34 => "0000",
		35 => "0000",
		36 => "1000",
		37 => "0000",
		38 => "0000",
		39 => "0000",
		40 => "1000",
		41 => "0000",
		42 => "0000",
		43 => "0000",
		44 => "0000",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 13
constant routing_table_bits_13: t_tata_long := (
	-- local
		0 => "0000",
		1 => "1000",
		2 => "0100",
		3 => "0000",
		4 => "0010",
		5 => "1000",
		6 => "0100",
		7 => "0000",
		8 => "0010",
		9 => "1000",
		10 => "0100",
		11 => "0000",
		12 => "0010",
		13 => "0000",
		14 => "0100",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0000",
		18 => "0100",
		19 => "0000",
		20 => "0010",
		21 => "0000",
		22 => "0100",
		23 => "0000",
		24 => "0010",
		25 => "0000",
		26 => "0100",
		27 => "0000",
		28 => "0010",
		29 => "0000",
		30 => "0100",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "1000",
		34 => "0000",
		35 => "0000",
		36 => "0010",
		37 => "1000",
		38 => "0000",
		39 => "0000",
		40 => "0010",
		41 => "1000",
		42 => "0000",
		43 => "0000",
		44 => "0010",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "1000",
		50 => "0100",
		51 => "0000",
		52 => "0000",
		53 => "1000",
		54 => "0100",
		55 => "0000",
		56 => "0000",
		57 => "1000",
		58 => "0100",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0100",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 14
constant routing_table_bits_14: t_tata_long := (
	-- local
		0 => "0000",
		1 => "0010",
		2 => "1000",
		3 => "0000",
		4 => "0010",
		5 => "0010",
		6 => "1000",
		7 => "0000",
		8 => "0010",
		9 => "0010",
		10 => "1000",
		11 => "0000",
		12 => "0010",
		13 => "0010",
		14 => "0000",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0010",
		18 => "0000",
		19 => "0000",
		20 => "0010",
		21 => "0010",
		22 => "0000",
		23 => "0000",
		24 => "0010",
		25 => "0010",
		26 => "0000",
		27 => "0000",
		28 => "0010",
		29 => "0010",
		30 => "0000",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "0000",
		34 => "0000",
		35 => "0000",
		36 => "0000",
		37 => "0000",
		38 => "0000",
		39 => "0000",
		40 => "0000",
		41 => "0000",
		42 => "0000",
		43 => "0000",
		44 => "0000",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "1000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "1000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "1000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );
-- Node 15
constant routing_table_bits_15: t_tata_long := (
	-- local
		0 => "1000",
		1 => "0000",
		2 => "0000",
		3 => "0000",
		4 => "0000",
		5 => "0000",
		6 => "0000",
		7 => "0000",
		8 => "0000",
		9 => "0000",
		10 => "0000",
		11 => "0000",
		12 => "0000",
		13 => "0000",
		14 => "0000",
		15 => "0000",
	-- north
		16 => "0000",
		17 => "0000",
		18 => "0000",
		19 => "0000",
		20 => "0000",
		21 => "0000",
		22 => "0000",
		23 => "0000",
		24 => "0000",
		25 => "0000",
		26 => "0000",
		27 => "0000",
		28 => "0000",
		29 => "0000",
		30 => "0000",
		31 => "0000",
	-- east
		32 => "0000",
		33 => "0000",
		34 => "0000",
		35 => "0000",
		36 => "0000",
		37 => "0000",
		38 => "0000",
		39 => "0000",
		40 => "0000",
		41 => "0000",
		42 => "0000",
		43 => "0000",
		44 => "0000",
		45 => "0000",
		46 => "0000",
		47 => "0000",
	-- west
		48 => "0000",
		49 => "0000",
		50 => "0000",
		51 => "0000",
		52 => "0000",
		53 => "0000",
		54 => "0000",
		55 => "0000",
		56 => "0000",
		57 => "0000",
		58 => "0000",
		59 => "0000",
		60 => "0000",
		61 => "0000",
		62 => "0000",
		63 => "0000",
	-- south
		64 => "0000",
		65 => "0000",
		66 => "0000",
		67 => "0000",
		68 => "0000",
		69 => "0000",
		70 => "0000",
		71 => "0000",
		72 => "0000",
		73 => "0000",
		74 => "0000",
		75 => "0000",
		76 => "0000",
		77 => "0000",
		78 => "0000",
		79 => "0000"
 );


--        organizaiton of the network:
--     x --------------->
--  y         ----       ----       ----       ----
--  |        | 0  | --- | 1  | --- | 2  | --- | 3  |
--  |         ----       ----       ----       ----
--  |          |          |          |          |
--  |         ----       ----       ----       ----
--  |        | 4  | --- | 5  | --- | 6  | --- | 7  |
--  |         ----       ----       ----       ----
--  |          |          |          |          |
--  |         ----       ----       ----       ----
--  |        | 8  | --- | 9  | --- | 10 | --- | 11 |
--  |         ----       ----       ----       ----
--  |          |          |          |          |
--  |         ----       ----       ----       ----
--  |        | 12 | --- | 13 | --- | 14 | --- | 15 |
--  v         ----       ----       ----       ----
--                                               
begin


-- instantiating the routers
R_0: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>0, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_0 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_0 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_0 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_0 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_0 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_0, RX_E_0, RX_W_0, RX_S_0, RX_L_0,
	credit_in_N_0, credit_in_E_0, credit_in_W_0, credit_in_S_0, credit_in_L_0,
	valid_in_N_0, valid_in_E_0, valid_in_W_0, valid_in_S_0, valid_in_L_0,
	valid_out_N_0, valid_out_E_0, valid_out_W_0, valid_out_S_0, valid_out_L_0,
	credit_out_N_0, credit_out_E_0, credit_out_W_0, credit_out_S_0, credit_out_L_0,
	TX_N_0, TX_E_0, TX_W_0, TX_S_0, TX_L_0); 

R_1: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>1, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_1 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_1 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_1 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_1 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_1 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_1, RX_E_1, RX_W_1, RX_S_1, RX_L_1,
	credit_in_N_1, credit_in_E_1, credit_in_W_1, credit_in_S_1, credit_in_L_1,
	valid_in_N_1, valid_in_E_1, valid_in_W_1, valid_in_S_1, valid_in_L_1,
	valid_out_N_1, valid_out_E_1, valid_out_W_1, valid_out_S_1, valid_out_L_1,
	credit_out_N_1, credit_out_E_1, credit_out_W_1, credit_out_S_1, credit_out_L_1,
	TX_N_1, TX_E_1, TX_W_1, TX_S_1, TX_L_1); 

R_2: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>2, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_2 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_2 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_2 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_2 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_2 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_2, RX_E_2, RX_W_2, RX_S_2, RX_L_2,
	credit_in_N_2, credit_in_E_2, credit_in_W_2, credit_in_S_2, credit_in_L_2,
	valid_in_N_2, valid_in_E_2, valid_in_W_2, valid_in_S_2, valid_in_L_2,
	valid_out_N_2, valid_out_E_2, valid_out_W_2, valid_out_S_2, valid_out_L_2,
	credit_out_N_2, credit_out_E_2, credit_out_W_2, credit_out_S_2, credit_out_L_2,
	TX_N_2, TX_E_2, TX_W_2, TX_S_2, TX_L_2); 

R_3: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>3, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_3 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_3 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_3 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_3 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_3 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_3, RX_E_3, RX_W_3, RX_S_3, RX_L_3,
	credit_in_N_3, credit_in_E_3, credit_in_W_3, credit_in_S_3, credit_in_L_3,
	valid_in_N_3, valid_in_E_3, valid_in_W_3, valid_in_S_3, valid_in_L_3,
	valid_out_N_3, valid_out_E_3, valid_out_W_3, valid_out_S_3, valid_out_L_3,
	credit_out_N_3, credit_out_E_3, credit_out_W_3, credit_out_S_3, credit_out_L_3,
	TX_N_3, TX_E_3, TX_W_3, TX_S_3, TX_L_3); 

R_4: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>4, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_4 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_4 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_4 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_4 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_4 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_4, RX_E_4, RX_W_4, RX_S_4, RX_L_4,
	credit_in_N_4, credit_in_E_4, credit_in_W_4, credit_in_S_4, credit_in_L_4,
	valid_in_N_4, valid_in_E_4, valid_in_W_4, valid_in_S_4, valid_in_L_4,
	valid_out_N_4, valid_out_E_4, valid_out_W_4, valid_out_S_4, valid_out_L_4,
	credit_out_N_4, credit_out_E_4, credit_out_W_4, credit_out_S_4, credit_out_L_4,
	TX_N_4, TX_E_4, TX_W_4, TX_S_4, TX_L_4); 

R_5: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>5, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_5 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_5 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_5 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_5 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_5 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_5, RX_E_5, RX_W_5, RX_S_5, RX_L_5,
	credit_in_N_5, credit_in_E_5, credit_in_W_5, credit_in_S_5, credit_in_L_5,
	valid_in_N_5, valid_in_E_5, valid_in_W_5, valid_in_S_5, valid_in_L_5,
	valid_out_N_5, valid_out_E_5, valid_out_W_5, valid_out_S_5, valid_out_L_5,
	credit_out_N_5, credit_out_E_5, credit_out_W_5, credit_out_S_5, credit_out_L_5,
	TX_N_5, TX_E_5, TX_W_5, TX_S_5, TX_L_5); 

R_6: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>6, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_6 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_6 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_6 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_6 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_6 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_6, RX_E_6, RX_W_6, RX_S_6, RX_L_6,
	credit_in_N_6, credit_in_E_6, credit_in_W_6, credit_in_S_6, credit_in_L_6,
	valid_in_N_6, valid_in_E_6, valid_in_W_6, valid_in_S_6, valid_in_L_6,
	valid_out_N_6, valid_out_E_6, valid_out_W_6, valid_out_S_6, valid_out_L_6,
	credit_out_N_6, credit_out_E_6, credit_out_W_6, credit_out_S_6, credit_out_L_6,
	TX_N_6, TX_E_6, TX_W_6, TX_S_6, TX_L_6); 

R_7: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>7, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_7 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_7 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_7 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_7 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_7 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_7, RX_E_7, RX_W_7, RX_S_7, RX_L_7,
	credit_in_N_7, credit_in_E_7, credit_in_W_7, credit_in_S_7, credit_in_L_7,
	valid_in_N_7, valid_in_E_7, valid_in_W_7, valid_in_S_7, valid_in_L_7,
	valid_out_N_7, valid_out_E_7, valid_out_W_7, valid_out_S_7, valid_out_L_7,
	credit_out_N_7, credit_out_E_7, credit_out_W_7, credit_out_S_7, credit_out_L_7,
	TX_N_7, TX_E_7, TX_W_7, TX_S_7, TX_L_7); 

R_8: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>8, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_8 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_8 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_8 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_8 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_8 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_8, RX_E_8, RX_W_8, RX_S_8, RX_L_8,
	credit_in_N_8, credit_in_E_8, credit_in_W_8, credit_in_S_8, credit_in_L_8,
	valid_in_N_8, valid_in_E_8, valid_in_W_8, valid_in_S_8, valid_in_L_8,
	valid_out_N_8, valid_out_E_8, valid_out_W_8, valid_out_S_8, valid_out_L_8,
	credit_out_N_8, credit_out_E_8, credit_out_W_8, credit_out_S_8, credit_out_L_8,
	TX_N_8, TX_E_8, TX_W_8, TX_S_8, TX_L_8); 

R_9: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>9, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_9 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_9 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_9 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_9 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_9 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_9, RX_E_9, RX_W_9, RX_S_9, RX_L_9,
	credit_in_N_9, credit_in_E_9, credit_in_W_9, credit_in_S_9, credit_in_L_9,
	valid_in_N_9, valid_in_E_9, valid_in_W_9, valid_in_S_9, valid_in_L_9,
	valid_out_N_9, valid_out_E_9, valid_out_W_9, valid_out_S_9, valid_out_L_9,
	credit_out_N_9, credit_out_E_9, credit_out_W_9, credit_out_S_9, credit_out_L_9,
	TX_N_9, TX_E_9, TX_W_9, TX_S_9, TX_L_9); 

R_10: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>10, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_10 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_10 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_10 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_10 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_10 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_10, RX_E_10, RX_W_10, RX_S_10, RX_L_10,
	credit_in_N_10, credit_in_E_10, credit_in_W_10, credit_in_S_10, credit_in_L_10,
	valid_in_N_10, valid_in_E_10, valid_in_W_10, valid_in_S_10, valid_in_L_10,
	valid_out_N_10, valid_out_E_10, valid_out_W_10, valid_out_S_10, valid_out_L_10,
	credit_out_N_10, credit_out_E_10, credit_out_W_10, credit_out_S_10, credit_out_L_10,
	TX_N_10, TX_E_10, TX_W_10, TX_S_10, TX_L_10); 

R_11: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>11, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_11 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_11 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_11 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_11 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_11 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_11, RX_E_11, RX_W_11, RX_S_11, RX_L_11,
	credit_in_N_11, credit_in_E_11, credit_in_W_11, credit_in_S_11, credit_in_L_11,
	valid_in_N_11, valid_in_E_11, valid_in_W_11, valid_in_S_11, valid_in_L_11,
	valid_out_N_11, valid_out_E_11, valid_out_W_11, valid_out_S_11, valid_out_L_11,
	credit_out_N_11, credit_out_E_11, credit_out_W_11, credit_out_S_11, credit_out_L_11,
	TX_N_11, TX_E_11, TX_W_11, TX_S_11, TX_L_11); 

R_12: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>12, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_12 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_12 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_12 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_12 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_12 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_12, RX_E_12, RX_W_12, RX_S_12, RX_L_12,
	credit_in_N_12, credit_in_E_12, credit_in_W_12, credit_in_S_12, credit_in_L_12,
	valid_in_N_12, valid_in_E_12, valid_in_W_12, valid_in_S_12, valid_in_L_12,
	valid_out_N_12, valid_out_E_12, valid_out_W_12, valid_out_S_12, valid_out_L_12,
	credit_out_N_12, credit_out_E_12, credit_out_W_12, credit_out_S_12, credit_out_L_12,
	TX_N_12, TX_E_12, TX_W_12, TX_S_12, TX_L_12); 

R_13: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>13, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_13 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_13 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_13 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_13 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_13 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_13, RX_E_13, RX_W_13, RX_S_13, RX_L_13,
	credit_in_N_13, credit_in_E_13, credit_in_W_13, credit_in_S_13, credit_in_L_13,
	valid_in_N_13, valid_in_E_13, valid_in_W_13, valid_in_S_13, valid_in_L_13,
	valid_out_N_13, valid_out_E_13, valid_out_W_13, valid_out_S_13, valid_out_L_13,
	credit_out_N_13, credit_out_E_13, credit_out_W_13, credit_out_S_13, credit_out_L_13,
	TX_N_13, TX_E_13, TX_W_13, TX_S_13, TX_L_13); 

R_14: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>14, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_14 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_14 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_14 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_14 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_14 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_14, RX_E_14, RX_W_14, RX_S_14, RX_L_14,
	credit_in_N_14, credit_in_E_14, credit_in_W_14, credit_in_S_14, credit_in_L_14,
	valid_in_N_14, valid_in_E_14, valid_in_W_14, valid_in_S_14, valid_in_L_14,
	valid_out_N_14, valid_out_E_14, valid_out_W_14, valid_out_S_14, valid_out_L_14,
	credit_out_N_14, credit_out_E_14, credit_out_W_14, credit_out_S_14, credit_out_L_14,
	TX_N_14, TX_E_14, TX_W_14, TX_S_14, TX_L_14); 

R_15: router_credit_based generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>15, NoC_size=>4, 
	routing_table_bits_local => t_tata (routing_table_bits_15 (0 to 15)), routing_table_bits_north => t_tata (routing_table_bits_15 (16 to 31)), 
	routing_table_bits_east => t_tata (routing_table_bits_15 (32 to 47)), routing_table_bits_west => t_tata (routing_table_bits_15 (48 to 63)), 
	routing_table_bits_south => t_tata (routing_table_bits_15 (64 to 79)))
PORT MAP (reset, clk, 
	RX_N_15, RX_E_15, RX_W_15, RX_S_15, RX_L_15,
	credit_in_N_15, credit_in_E_15, credit_in_W_15, credit_in_S_15, credit_in_L_15,
	valid_in_N_15, valid_in_E_15, valid_in_W_15, valid_in_S_15, valid_in_L_15,
	valid_out_N_15, valid_out_E_15, valid_out_W_15, valid_out_S_15, valid_out_L_15,
	credit_out_N_15, credit_out_E_15, credit_out_W_15, credit_out_S_15, credit_out_L_15,
	TX_N_15, TX_E_15, TX_W_15, TX_S_15, TX_L_15); 


---------------------------------------------------------------
-- binding the routers together
-- vertical ins/outs
-- connecting router: 0 to router: 4 and vice versa
RX_N_4<= TX_S_0;
RX_S_0<= TX_N_4;
-------------------
-- connecting router: 1 to router: 5 and vice versa
RX_N_5<= TX_S_1;
RX_S_1<= TX_N_5;
-------------------
-- connecting router: 2 to router: 6 and vice versa
RX_N_6<= TX_S_2;
RX_S_2<= TX_N_6;
-------------------
-- connecting router: 3 to router: 7 and vice versa
RX_N_7<= TX_S_3;
RX_S_3<= TX_N_7;
-------------------
-- connecting router: 4 to router: 8 and vice versa
RX_N_8<= TX_S_4;
RX_S_4<= TX_N_8;
-------------------
-- connecting router: 5 to router: 9 and vice versa
RX_N_9<= TX_S_5;
RX_S_5<= TX_N_9;
-------------------
-- connecting router: 6 to router: 10 and vice versa
RX_N_10<= TX_S_6;
RX_S_6<= TX_N_10;
-------------------
-- connecting router: 7 to router: 11 and vice versa
RX_N_11<= TX_S_7;
RX_S_7<= TX_N_11;
-------------------
-- connecting router: 8 to router: 12 and vice versa
RX_N_12<= TX_S_8;
RX_S_8<= TX_N_12;
-------------------
-- connecting router: 9 to router: 13 and vice versa
RX_N_13<= TX_S_9;
RX_S_9<= TX_N_13;
-------------------
-- connecting router: 10 to router: 14 and vice versa
RX_N_14<= TX_S_10;
RX_S_10<= TX_N_14;
-------------------
-- connecting router: 11 to router: 15 and vice versa
RX_N_15<= TX_S_11;
RX_S_11<= TX_N_15;
-------------------

-- horizontal ins/outs
-- connecting router: 0 to router: 1 and vice versa
RX_E_0 <= TX_W_1;
RX_W_1 <= TX_E_0;
-------------------
-- connecting router: 1 to router: 2 and vice versa
RX_E_1 <= TX_W_2;
RX_W_2 <= TX_E_1;
-------------------
-- connecting router: 2 to router: 3 and vice versa
RX_E_2 <= TX_W_3;
RX_W_3 <= TX_E_2;
-------------------
-- connecting router: 4 to router: 5 and vice versa
RX_E_4 <= TX_W_5;
RX_W_5 <= TX_E_4;
-------------------
-- connecting router: 5 to router: 6 and vice versa
RX_E_5 <= TX_W_6;
RX_W_6 <= TX_E_5;
-------------------
-- connecting router: 6 to router: 7 and vice versa
RX_E_6 <= TX_W_7;
RX_W_7 <= TX_E_6;
-------------------
-- connecting router: 8 to router: 9 and vice versa
RX_E_8 <= TX_W_9;
RX_W_9 <= TX_E_8;
-------------------
-- connecting router: 9 to router: 10 and vice versa
RX_E_9 <= TX_W_10;
RX_W_10 <= TX_E_9;
-------------------
-- connecting router: 10 to router: 11 and vice versa
RX_E_10 <= TX_W_11;
RX_W_11 <= TX_E_10;
-------------------
-- connecting router: 12 to router: 13 and vice versa
RX_E_12 <= TX_W_13;
RX_W_13 <= TX_E_12;
-------------------
-- connecting router: 13 to router: 14 and vice versa
RX_E_13 <= TX_W_14;
RX_W_14 <= TX_E_13;
-------------------
-- connecting router: 14 to router: 15 and vice versa
RX_E_14 <= TX_W_15;
RX_W_15 <= TX_E_14;
-------------------
---------------------------------------------------------------
-- binding the routers together
-- connecting router: 0 to router: 4 and vice versa
valid_in_N_4 <= valid_out_S_0;
valid_in_S_0 <= valid_out_N_4;
credit_in_S_0 <= credit_out_N_4;
credit_in_N_4 <= credit_out_S_0;
-------------------
-- connecting router: 1 to router: 5 and vice versa
valid_in_N_5 <= valid_out_S_1;
valid_in_S_1 <= valid_out_N_5;
credit_in_S_1 <= credit_out_N_5;
credit_in_N_5 <= credit_out_S_1;
-------------------
-- connecting router: 2 to router: 6 and vice versa
valid_in_N_6 <= valid_out_S_2;
valid_in_S_2 <= valid_out_N_6;
credit_in_S_2 <= credit_out_N_6;
credit_in_N_6 <= credit_out_S_2;
-------------------
-- connecting router: 3 to router: 7 and vice versa
valid_in_N_7 <= valid_out_S_3;
valid_in_S_3 <= valid_out_N_7;
credit_in_S_3 <= credit_out_N_7;
credit_in_N_7 <= credit_out_S_3;
-------------------
-- connecting router: 4 to router: 8 and vice versa
valid_in_N_8 <= valid_out_S_4;
valid_in_S_4 <= valid_out_N_8;
credit_in_S_4 <= credit_out_N_8;
credit_in_N_8 <= credit_out_S_4;
-------------------
-- connecting router: 5 to router: 9 and vice versa
valid_in_N_9 <= valid_out_S_5;
valid_in_S_5 <= valid_out_N_9;
credit_in_S_5 <= credit_out_N_9;
credit_in_N_9 <= credit_out_S_5;
-------------------
-- connecting router: 6 to router: 10 and vice versa
valid_in_N_10 <= valid_out_S_6;
valid_in_S_6 <= valid_out_N_10;
credit_in_S_6 <= credit_out_N_10;
credit_in_N_10 <= credit_out_S_6;
-------------------
-- connecting router: 7 to router: 11 and vice versa
valid_in_N_11 <= valid_out_S_7;
valid_in_S_7 <= valid_out_N_11;
credit_in_S_7 <= credit_out_N_11;
credit_in_N_11 <= credit_out_S_7;
-------------------
-- connecting router: 8 to router: 12 and vice versa
valid_in_N_12 <= valid_out_S_8;
valid_in_S_8 <= valid_out_N_12;
credit_in_S_8 <= credit_out_N_12;
credit_in_N_12 <= credit_out_S_8;
-------------------
-- connecting router: 9 to router: 13 and vice versa
valid_in_N_13 <= valid_out_S_9;
valid_in_S_9 <= valid_out_N_13;
credit_in_S_9 <= credit_out_N_13;
credit_in_N_13 <= credit_out_S_9;
-------------------
-- connecting router: 10 to router: 14 and vice versa
valid_in_N_14 <= valid_out_S_10;
valid_in_S_10 <= valid_out_N_14;
credit_in_S_10 <= credit_out_N_14;
credit_in_N_14 <= credit_out_S_10;
-------------------
-- connecting router: 11 to router: 15 and vice versa
valid_in_N_15 <= valid_out_S_11;
valid_in_S_11 <= valid_out_N_15;
credit_in_S_11 <= credit_out_N_15;
credit_in_N_15 <= credit_out_S_11;
-------------------

-- connecting router: 0 to router: 1 and vice versa
valid_in_E_0 <= valid_out_W_1;
valid_in_W_1 <= valid_out_E_0;
credit_in_W_1 <= credit_out_E_0;
credit_in_E_0 <= credit_out_W_1;
-------------------
-- connecting router: 1 to router: 2 and vice versa
valid_in_E_1 <= valid_out_W_2;
valid_in_W_2 <= valid_out_E_1;
credit_in_W_2 <= credit_out_E_1;
credit_in_E_1 <= credit_out_W_2;
-------------------
-- connecting router: 2 to router: 3 and vice versa
valid_in_E_2 <= valid_out_W_3;
valid_in_W_3 <= valid_out_E_2;
credit_in_W_3 <= credit_out_E_2;
credit_in_E_2 <= credit_out_W_3;
-------------------
-- connecting router: 4 to router: 5 and vice versa
valid_in_E_4 <= valid_out_W_5;
valid_in_W_5 <= valid_out_E_4;
credit_in_W_5 <= credit_out_E_4;
credit_in_E_4 <= credit_out_W_5;
-------------------
-- connecting router: 5 to router: 6 and vice versa
valid_in_E_5 <= valid_out_W_6;
valid_in_W_6 <= valid_out_E_5;
credit_in_W_6 <= credit_out_E_5;
credit_in_E_5 <= credit_out_W_6;
-------------------
-- connecting router: 6 to router: 7 and vice versa
valid_in_E_6 <= valid_out_W_7;
valid_in_W_7 <= valid_out_E_6;
credit_in_W_7 <= credit_out_E_6;
credit_in_E_6 <= credit_out_W_7;
-------------------
-- connecting router: 8 to router: 9 and vice versa
valid_in_E_8 <= valid_out_W_9;
valid_in_W_9 <= valid_out_E_8;
credit_in_W_9 <= credit_out_E_8;
credit_in_E_8 <= credit_out_W_9;
-------------------
-- connecting router: 9 to router: 10 and vice versa
valid_in_E_9 <= valid_out_W_10;
valid_in_W_10 <= valid_out_E_9;
credit_in_W_10 <= credit_out_E_9;
credit_in_E_9 <= credit_out_W_10;
-------------------
-- connecting router: 10 to router: 11 and vice versa
valid_in_E_10 <= valid_out_W_11;
valid_in_W_11 <= valid_out_E_10;
credit_in_W_11 <= credit_out_E_10;
credit_in_E_10 <= credit_out_W_11;
-------------------
-- connecting router: 12 to router: 13 and vice versa
valid_in_E_12 <= valid_out_W_13;
valid_in_W_13 <= valid_out_E_12;
credit_in_W_13 <= credit_out_E_12;
credit_in_E_12 <= credit_out_W_13;
-------------------
-- connecting router: 13 to router: 14 and vice versa
valid_in_E_13 <= valid_out_W_14;
valid_in_W_14 <= valid_out_E_13;
credit_in_W_14 <= credit_out_E_13;
credit_in_E_13 <= credit_out_W_14;
-------------------
-- connecting router: 14 to router: 15 and vice versa
valid_in_E_14 <= valid_out_W_15;
valid_in_W_15 <= valid_out_E_14;
credit_in_W_15 <= credit_out_E_14;
credit_in_E_14 <= credit_out_W_15;
-------------------
end;
