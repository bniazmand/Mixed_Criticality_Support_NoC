--Copyright (C) 2016 Siavoosh Payandeh Azad

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.all;
 use ieee.math_real.all;
 use std.textio.all;
 use ieee.std_logic_misc.all;

package type_def_pack is

   type t_tata IS ARRAY(0 to 15) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
   type t_tata_long IS ARRAY(0 to 79) OF STD_LOGIC_VECTOR(3 DOWNTO 0);

  -- Node 0
   constant routing_table_bits_0: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "0000",
   		5 => "0000",
   		6 => "0000",
   		7 => "0000",
   		8 => "0000",
   		9 => "0000",
   		10 => "0000",
   		11 => "0000",
   		12 => "0000",
   		13 => "0000",
   		14 => "0000",
   		15 => "0100",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 1
   constant routing_table_bits_1: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0100",
   		3 => "0100",
   		4 => "0100",
   		5 => "0100",
   		6 => "0100",
   		7 => "0100",
   		8 => "0100",
   		9 => "0100",
   		10 => "0100",
   		11 => "0100",
   		12 => "0100",
   		13 => "0100",
   		14 => "0100",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0001",
   	-- south
   		64 => "0010",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 2
   constant routing_table_bits_2: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0010",
   		2 => "0000",
   		3 => "0100",
   		4 => "0101",
   		5 => "0101",
   		6 => "0101",
   		7 => "0101",
   		8 => "0101",
   		9 => "0101",
   		10 => "0101",
   		11 => "0101",
   		12 => "0101",
   		13 => "0101",
   		14 => "0101",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0010",
   		34 => "0000",
   		35 => "0000",
   		36 => "0001",
   		37 => "0001",
   		38 => "0001",
   		39 => "0001",
   		40 => "0001",
   		41 => "0001",
   		42 => "0001",
   		43 => "0001",
   		44 => "0001",
   		45 => "0001",
   		46 => "0001",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0100",
   		52 => "0101",
   		53 => "0101",
   		54 => "0101",
   		55 => "0101",
   		56 => "0101",
   		57 => "0101",
   		58 => "0101",
   		59 => "0101",
   		60 => "0101",
   		61 => "0101",
   		62 => "0101",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0010",
   		66 => "0000",
   		67 => "0100",
   		68 => "0100",
   		69 => "0100",
   		70 => "0100",
   		71 => "0100",
   		72 => "0100",
   		73 => "0100",
   		74 => "0100",
   		75 => "0100",
   		76 => "0100",
   		77 => "0100",
   		78 => "0100",
   		79 => "0000"
    );
   -- Node 3
   constant routing_table_bits_3: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0010",
   		2 => "0010",
   		3 => "0000",
   		4 => "0011",
   		5 => "0011",
   		6 => "0011",
   		7 => "0011",
   		8 => "0011",
   		9 => "0011",
   		10 => "0011",
   		11 => "0011",
   		12 => "0011",
   		13 => "0011",
   		14 => "0011",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0001",
   		53 => "0001",
   		54 => "0001",
   		55 => "0001",
   		56 => "0001",
   		57 => "0001",
   		58 => "0001",
   		59 => "0001",
   		60 => "0001",
   		61 => "0001",
   		62 => "0001",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0010",
   		66 => "0010",
   		67 => "0000",
   		68 => "0010",
   		69 => "0010",
   		70 => "0010",
   		71 => "0010",
   		72 => "0010",
   		73 => "0010",
   		74 => "0010",
   		75 => "0010",
   		76 => "0010",
   		77 => "0010",
   		78 => "0010",
   		79 => "0000"
    );
   -- Node 4
   constant routing_table_bits_4: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "0000",
   		5 => "0100",
   		6 => "0100",
   		7 => "0100",
   		8 => "0001",
   		9 => "0001",
   		10 => "0100",
   		11 => "0100",
   		12 => "0001",
   		13 => "0001",
   		14 => "0001",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0001",
   		41 => "0001",
   		42 => "0000",
   		43 => "0000",
   		44 => "0001",
   		45 => "0001",
   		46 => "0001",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0100",
   		70 => "0100",
   		71 => "0100",
   		72 => "0000",
   		73 => "0000",
   		74 => "0100",
   		75 => "0100",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 5
   constant routing_table_bits_5: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "0010",
   		5 => "0000",
   		6 => "0100",
   		7 => "0100",
   		8 => "0010",
   		9 => "0010",
   		10 => "0100",
   		11 => "0100",
   		12 => "0010",
   		13 => "0010",
   		14 => "0010",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0001",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0010",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0010",
   		41 => "0010",
   		42 => "0000",
   		43 => "0000",
   		44 => "0010",
   		45 => "0010",
   		46 => "0010",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0100",
   		55 => "0100",
   		56 => "0000",
   		57 => "0000",
   		58 => "0100",
   		59 => "0100",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "1000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 6
   constant routing_table_bits_6: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "1000",
   		2 => "1000",
   		3 => "1000",
   		4 => "1010",
   		5 => "1010",
   		6 => "0000",
   		7 => "1100",
   		8 => "1010",
   		9 => "1010",
   		10 => "0101",
   		11 => "0101",
   		12 => "1010",
   		13 => "1010",
   		14 => "1010",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0010",
   		21 => "0010",
   		22 => "0000",
   		23 => "0100",
   		24 => "0010",
   		25 => "0010",
   		26 => "0101",
   		27 => "0101",
   		28 => "0010",
   		29 => "0010",
   		30 => "0010",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0010",
   		37 => "0010",
   		38 => "0000",
   		39 => "0000",
   		40 => "0010",
   		41 => "0010",
   		42 => "0001",
   		43 => "0001",
   		44 => "0010",
   		45 => "0010",
   		46 => "0010",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0100",
   		56 => "0000",
   		57 => "0000",
   		58 => "0101",
   		59 => "0101",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "1000",
   		66 => "1000",
   		67 => "1000",
   		68 => "1010",
   		69 => "1010",
   		70 => "0000",
   		71 => "1100",
   		72 => "1010",
   		73 => "1010",
   		74 => "1100",
   		75 => "1100",
   		76 => "1010",
   		77 => "1010",
   		78 => "1010",
   		79 => "0000"
    );
   -- Node 7
   constant routing_table_bits_7: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "1000",
   		2 => "1000",
   		3 => "1000",
   		4 => "1010",
   		5 => "1010",
   		6 => "1010",
   		7 => "0000",
   		8 => "1010",
   		9 => "1010",
   		10 => "0011",
   		11 => "0011",
   		12 => "1010",
   		13 => "1010",
   		14 => "1010",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0010",
   		21 => "0010",
   		22 => "0010",
   		23 => "0000",
   		24 => "0010",
   		25 => "0010",
   		26 => "0011",
   		27 => "0011",
   		28 => "0010",
   		29 => "0010",
   		30 => "0010",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0001",
   		59 => "0001",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "1000",
   		66 => "1000",
   		67 => "1000",
   		68 => "1010",
   		69 => "1010",
   		70 => "1010",
   		71 => "0000",
   		72 => "1010",
   		73 => "1010",
   		74 => "1010",
   		75 => "1010",
   		76 => "1010",
   		77 => "1010",
   		78 => "1010",
   		79 => "0000"
    );
   -- Node 8
   constant routing_table_bits_8: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "1000",
   		5 => "1000",
   		6 => "1000",
   		7 => "1000",
   		8 => "0000",
   		9 => "0100",
   		10 => "1000",
   		11 => "1000",
   		12 => "0101",
   		13 => "0101",
   		14 => "0101",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0100",
   		26 => "0000",
   		27 => "0000",
   		28 => "0101",
   		29 => "0101",
   		30 => "0101",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0001",
   		45 => "0001",
   		46 => "0001",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "1000",
   		69 => "1000",
   		70 => "1000",
   		71 => "1000",
   		72 => "0000",
   		73 => "0100",
   		74 => "1000",
   		75 => "1000",
   		76 => "0100",
   		77 => "0100",
   		78 => "0100",
   		79 => "0000"
    );
   -- Node 9
   constant routing_table_bits_9: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "0000",
   		5 => "0000",
   		6 => "0000",
   		7 => "0000",
   		8 => "0010",
   		9 => "0000",
   		10 => "0000",
   		11 => "0000",
   		12 => "0011",
   		13 => "0011",
   		14 => "0011",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0100",
   	-- east
   		32 => "1000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0001",
   		61 => "0001",
   		62 => "0001",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0010",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0010",
   		77 => "0010",
   		78 => "0010",
   		79 => "0000"
    );
   -- Node 10
   constant routing_table_bits_10: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "1000",
   		2 => "1000",
   		3 => "1000",
   		4 => "1000",
   		5 => "1000",
   		6 => "1000",
   		7 => "1000",
   		8 => "1000",
   		9 => "1000",
   		10 => "0000",
   		11 => "1100",
   		12 => "1000",
   		13 => "1000",
   		14 => "1000",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0100",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0001",
   	-- south
   		64 => "0010",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 11
   constant routing_table_bits_11: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "1000",
   		2 => "1000",
   		3 => "1000",
   		4 => "1000",
   		5 => "1000",
   		6 => "1000",
   		7 => "1000",
   		8 => "1000",
   		9 => "1000",
   		10 => "1010",
   		11 => "0000",
   		12 => "1000",
   		13 => "1000",
   		14 => "1000",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0010",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 12
   constant routing_table_bits_12: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "1000",
   		5 => "1000",
   		6 => "1000",
   		7 => "1000",
   		8 => "1000",
   		9 => "1000",
   		10 => "1000",
   		11 => "1000",
   		12 => "0000",
   		13 => "1100",
   		14 => "1100",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0100",
   		30 => "0100",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 13
   constant routing_table_bits_13: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "0000",
   		5 => "0000",
   		6 => "0000",
   		7 => "0000",
   		8 => "1000",
   		9 => "1000",
   		10 => "0000",
   		11 => "0000",
   		12 => "1010",
   		13 => "0000",
   		14 => "1100",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0010",
   		29 => "0000",
   		30 => "0100",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0010",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0100",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 14
   constant routing_table_bits_14: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "0000",
   		5 => "0000",
   		6 => "0000",
   		7 => "0000",
   		8 => "0000",
   		9 => "0000",
   		10 => "0000",
   		11 => "0000",
   		12 => "0010",
   		13 => "0010",
   		14 => "0000",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0100",
   	-- east
   		32 => "1000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 15
   constant routing_table_bits_15: t_tata_long := (
   	-- local
   		0 => "0010",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "0000",
   		5 => "0000",
   		6 => "0000",
   		7 => "0000",
   		8 => "0000",
   		9 => "0000",
   		10 => "0000",
   		11 => "0000",
   		12 => "0000",
   		13 => "0000",
   		14 => "0000",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );


 constant sel_N_R_0 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_0 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_0 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_0 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_1 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_1 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_1 : std_logic_vector(1 downto 0):=  "01";
 constant sel_S_R_1 : std_logic_vector(1 downto 0):=  "11";

 constant sel_N_R_2 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_2 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_2 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_2 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_3 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_3 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_3 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_3 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_4 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_4 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_4 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_4 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_5 : std_logic_vector(1 downto 0):=  "11";
 constant sel_E_R_5 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_5 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_5 : std_logic_vector(1 downto 0):=  "01";

 constant sel_N_R_6 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_6 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_6 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_6 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_7 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_7 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_7 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_7 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_8 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_8 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_8 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_8 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_9 : std_logic_vector(1 downto 0):=  "01";
 constant sel_E_R_9 : std_logic_vector(1 downto 0):=  "11";
 constant sel_W_R_9 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_9 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_10 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_10 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_10 : std_logic_vector(1 downto 0):=  "01";
 constant sel_S_R_10 : std_logic_vector(1 downto 0):=  "11";

 constant sel_N_R_11 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_11 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_11 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_11 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_12 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_12 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_12 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_12 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_13 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_13 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_13 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_13 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_14 : std_logic_vector(1 downto 0):=  "01";
 constant sel_E_R_14 : std_logic_vector(1 downto 0):=  "11";
 constant sel_W_R_14 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_14 : std_logic_vector(1 downto 0):=  "00";

 constant sel_N_R_15 : std_logic_vector(1 downto 0):=  "00";
 constant sel_E_R_15 : std_logic_vector(1 downto 0):=  "00";
 constant sel_W_R_15 : std_logic_vector(1 downto 0):=  "00";
 constant sel_S_R_15 : std_logic_vector(1 downto 0):=  "00";


end type_def_pack;
