--Copyright (C) 2016 Siavoosh Payandeh Azad

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.all;
 use ieee.math_real.all;
 use std.textio.all;
 use ieee.std_logic_misc.all;

package type_def_pack is

   type t_tata IS ARRAY(0 to 15) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
   type t_tata_long IS ARRAY(0 to 79) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
   -- Node 0
   constant routing_table_bits_0: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "0000",
   		5 => "0000",
   		6 => "0000",
   		7 => "0000",
   		8 => "0000",
   		9 => "0000",
   		10 => "0000",
   		11 => "0000",
   		12 => "0000",
   		13 => "0000",
   		14 => "0100",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 1
   constant routing_table_bits_1: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0000",
   		2 => "0001",
   		3 => "0001",
   		4 => "0001",
   		5 => "0001",
   		6 => "0001",
   		7 => "0001",
   		8 => "0001",
   		9 => "0001",
   		10 => "0001",
   		11 => "0001",
   		12 => "0001",
   		13 => "0001",
   		14 => "0000",
   		15 => "0001",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0010",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0100",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 2
   constant routing_table_bits_2: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0100",
   		2 => "0000",
   		3 => "0100",
   		4 => "0100",
   		5 => "0100",
   		6 => "0100",
   		7 => "0100",
   		8 => "0100",
   		9 => "0100",
   		10 => "0100",
   		11 => "0100",
   		12 => "0100",
   		13 => "0100",
   		14 => "0000",
   		15 => "0100",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0001",
   		63 => "0000",
   	-- south
   		64 => "0010",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 3
   constant routing_table_bits_3: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0001",
   		2 => "0010",
   		3 => "0000",
   		4 => "0001",
   		5 => "0001",
   		6 => "0001",
   		7 => "0001",
   		8 => "0001",
   		9 => "0001",
   		10 => "0001",
   		11 => "0001",
   		12 => "0001",
   		13 => "0001",
   		14 => "0000",
   		15 => "0001",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0001",
   		50 => "0000",
   		51 => "0000",
   		52 => "0001",
   		53 => "0001",
   		54 => "0001",
   		55 => "0001",
   		56 => "0001",
   		57 => "0001",
   		58 => "0001",
   		59 => "0001",
   		60 => "0001",
   		61 => "0001",
   		62 => "0000",
   		63 => "0001",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0010",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 4
   constant routing_table_bits_4: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0101",
   		2 => "0101",
   		3 => "0101",
   		4 => "0000",
   		5 => "0101",
   		6 => "0101",
   		7 => "0101",
   		8 => "0101",
   		9 => "0101",
   		10 => "0101",
   		11 => "0101",
   		12 => "0101",
   		13 => "0101",
   		14 => "0000",
   		15 => "0101",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 5
   constant routing_table_bits_5: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "1100",
   		2 => "0101",
   		3 => "0101",
   		4 => "0111",
   		5 => "0000",
   		6 => "0101",
   		7 => "0101",
   		8 => "0101",
   		9 => "0101",
   		10 => "0101",
   		11 => "0101",
   		12 => "0101",
   		13 => "0101",
   		14 => "0000",
   		15 => "0101",
   	-- north
   		16 => "0000",
   		17 => "0101",
   		18 => "0101",
   		19 => "0101",
   		20 => "0111",
   		21 => "0000",
   		22 => "0101",
   		23 => "0101",
   		24 => "0101",
   		25 => "0101",
   		26 => "0101",
   		27 => "0101",
   		28 => "0101",
   		29 => "0101",
   		30 => "0000",
   		31 => "0101",
   	-- east
   		32 => "0000",
   		33 => "1000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0010",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "1100",
   		50 => "0101",
   		51 => "0101",
   		52 => "0101",
   		53 => "0000",
   		54 => "0101",
   		55 => "0101",
   		56 => "0101",
   		57 => "0101",
   		58 => "0101",
   		59 => "0101",
   		60 => "0101",
   		61 => "0101",
   		62 => "0000",
   		63 => "0101",
   	-- south
   		64 => "0000",
   		65 => "1000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0010",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 6
   constant routing_table_bits_6: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0110",
   		2 => "0100",
   		3 => "0100",
   		4 => "0110",
   		5 => "0110",
   		6 => "0000",
   		7 => "0100",
   		8 => "0100",
   		9 => "0100",
   		10 => "0100",
   		11 => "0100",
   		12 => "0100",
   		13 => "0100",
   		14 => "0000",
   		15 => "0100",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0001",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0010",
   		34 => "0000",
   		35 => "0000",
   		36 => "0010",
   		37 => "0010",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0100",
   		50 => "0100",
   		51 => "0100",
   		52 => "0100",
   		53 => "0100",
   		54 => "0000",
   		55 => "0100",
   		56 => "0100",
   		57 => "0100",
   		58 => "0100",
   		59 => "0100",
   		60 => "0100",
   		61 => "0100",
   		62 => "0000",
   		63 => "0100",
   	-- south
   		64 => "1000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 7
   constant routing_table_bits_7: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0011",
   		2 => "1000",
   		3 => "1000",
   		4 => "0011",
   		5 => "0011",
   		6 => "0010",
   		7 => "0000",
   		8 => "0001",
   		9 => "0001",
   		10 => "0001",
   		11 => "0001",
   		12 => "0001",
   		13 => "0001",
   		14 => "0000",
   		15 => "0001",
   	-- north
   		16 => "0000",
   		17 => "0011",
   		18 => "0000",
   		19 => "0000",
   		20 => "0011",
   		21 => "0011",
   		22 => "0010",
   		23 => "0000",
   		24 => "0001",
   		25 => "0001",
   		26 => "0001",
   		27 => "0001",
   		28 => "0001",
   		29 => "0001",
   		30 => "0000",
   		31 => "0001",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0001",
   		50 => "1000",
   		51 => "1000",
   		52 => "0001",
   		53 => "0001",
   		54 => "0000",
   		55 => "0000",
   		56 => "0001",
   		57 => "0001",
   		58 => "0001",
   		59 => "0001",
   		60 => "0001",
   		61 => "0001",
   		62 => "0000",
   		63 => "0001",
   	-- south
   		64 => "0000",
   		65 => "0010",
   		66 => "1000",
   		67 => "1000",
   		68 => "0010",
   		69 => "0010",
   		70 => "0010",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 8
   constant routing_table_bits_8: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0101",
   		2 => "0101",
   		3 => "0101",
   		4 => "1100",
   		5 => "0101",
   		6 => "0101",
   		7 => "0101",
   		8 => "0000",
   		9 => "0101",
   		10 => "0101",
   		11 => "0101",
   		12 => "0101",
   		13 => "0101",
   		14 => "0000",
   		15 => "0101",
   	-- north
   		16 => "0000",
   		17 => "0101",
   		18 => "0101",
   		19 => "0101",
   		20 => "0101",
   		21 => "0101",
   		22 => "0101",
   		23 => "0101",
   		24 => "0000",
   		25 => "0101",
   		26 => "0101",
   		27 => "0101",
   		28 => "0101",
   		29 => "0101",
   		30 => "0000",
   		31 => "0101",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "1000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "1000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 9
   constant routing_table_bits_9: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0101",
   		2 => "0101",
   		3 => "0101",
   		4 => "0111",
   		5 => "0101",
   		6 => "0101",
   		7 => "0101",
   		8 => "0111",
   		9 => "0000",
   		10 => "0101",
   		11 => "0101",
   		12 => "0101",
   		13 => "0101",
   		14 => "0000",
   		15 => "0101",
   	-- north
   		16 => "0000",
   		17 => "0101",
   		18 => "0101",
   		19 => "0101",
   		20 => "0111",
   		21 => "0101",
   		22 => "0101",
   		23 => "0101",
   		24 => "0111",
   		25 => "0000",
   		26 => "0101",
   		27 => "0101",
   		28 => "0101",
   		29 => "0101",
   		30 => "0000",
   		31 => "0101",
   	-- east
   		32 => "0000",
   		33 => "1000",
   		34 => "0000",
   		35 => "0000",
   		36 => "1010",
   		37 => "1000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0010",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0101",
   		50 => "0101",
   		51 => "0101",
   		52 => "0101",
   		53 => "0101",
   		54 => "0101",
   		55 => "0101",
   		56 => "0101",
   		57 => "0000",
   		58 => "0101",
   		59 => "0101",
   		60 => "0101",
   		61 => "0101",
   		62 => "0000",
   		63 => "0101",
   	-- south
   		64 => "0000",
   		65 => "1000",
   		66 => "0000",
   		67 => "0000",
   		68 => "1010",
   		69 => "1000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0010",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 10
   constant routing_table_bits_10: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0110",
   		2 => "0100",
   		3 => "0100",
   		4 => "0110",
   		5 => "0110",
   		6 => "0100",
   		7 => "0100",
   		8 => "0110",
   		9 => "0110",
   		10 => "0000",
   		11 => "0100",
   		12 => "0100",
   		13 => "0100",
   		14 => "0000",
   		15 => "0100",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0001",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0010",
   		34 => "0000",
   		35 => "0000",
   		36 => "0010",
   		37 => "0010",
   		38 => "0000",
   		39 => "0000",
   		40 => "0010",
   		41 => "0010",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0100",
   		50 => "0100",
   		51 => "0100",
   		52 => "0100",
   		53 => "0100",
   		54 => "0100",
   		55 => "0100",
   		56 => "0100",
   		57 => "0100",
   		58 => "0000",
   		59 => "0100",
   		60 => "0100",
   		61 => "0100",
   		62 => "0000",
   		63 => "0100",
   	-- south
   		64 => "1000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 11
   constant routing_table_bits_11: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0011",
   		2 => "1000",
   		3 => "1000",
   		4 => "0011",
   		5 => "0011",
   		6 => "1000",
   		7 => "1000",
   		8 => "0011",
   		9 => "0011",
   		10 => "0010",
   		11 => "0000",
   		12 => "0001",
   		13 => "0001",
   		14 => "0000",
   		15 => "0001",
   	-- north
   		16 => "0000",
   		17 => "0011",
   		18 => "0000",
   		19 => "0000",
   		20 => "0011",
   		21 => "0011",
   		22 => "0000",
   		23 => "0000",
   		24 => "0011",
   		25 => "0011",
   		26 => "0010",
   		27 => "0000",
   		28 => "0001",
   		29 => "0001",
   		30 => "0000",
   		31 => "0001",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0001",
   		50 => "1000",
   		51 => "1000",
   		52 => "0001",
   		53 => "0001",
   		54 => "1000",
   		55 => "1000",
   		56 => "0001",
   		57 => "0001",
   		58 => "0000",
   		59 => "0000",
   		60 => "0001",
   		61 => "0001",
   		62 => "0000",
   		63 => "0001",
   	-- south
   		64 => "0000",
   		65 => "1010",
   		66 => "1000",
   		67 => "1000",
   		68 => "1010",
   		69 => "1010",
   		70 => "1000",
   		71 => "1000",
   		72 => "0010",
   		73 => "0010",
   		74 => "0010",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 12
   constant routing_table_bits_12: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "0100",
   		2 => "0100",
   		3 => "0100",
   		4 => "1100",
   		5 => "0100",
   		6 => "0100",
   		7 => "0100",
   		8 => "1100",
   		9 => "0100",
   		10 => "0100",
   		11 => "0100",
   		12 => "0000",
   		13 => "0100",
   		14 => "0000",
   		15 => "0100",
   	-- north
   		16 => "0000",
   		17 => "0100",
   		18 => "0100",
   		19 => "0100",
   		20 => "0100",
   		21 => "0100",
   		22 => "0100",
   		23 => "0100",
   		24 => "0100",
   		25 => "0100",
   		26 => "0100",
   		27 => "0100",
   		28 => "0000",
   		29 => "0100",
   		30 => "0000",
   		31 => "0100",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "1000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "1000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0000",
   		50 => "0000",
   		51 => "0000",
   		52 => "0000",
   		53 => "0000",
   		54 => "0000",
   		55 => "0000",
   		56 => "0000",
   		57 => "0000",
   		58 => "0000",
   		59 => "0000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 13
   constant routing_table_bits_13: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "1100",
   		2 => "0100",
   		3 => "0100",
   		4 => "1110",
   		5 => "1100",
   		6 => "0100",
   		7 => "0100",
   		8 => "1110",
   		9 => "1100",
   		10 => "0100",
   		11 => "0100",
   		12 => "0010",
   		13 => "0000",
   		14 => "0000",
   		15 => "0100",
   	-- north
   		16 => "0000",
   		17 => "0100",
   		18 => "0100",
   		19 => "0100",
   		20 => "0110",
   		21 => "0100",
   		22 => "0100",
   		23 => "0100",
   		24 => "0110",
   		25 => "0100",
   		26 => "0100",
   		27 => "0100",
   		28 => "0010",
   		29 => "0000",
   		30 => "0000",
   		31 => "0100",
   	-- east
   		32 => "0000",
   		33 => "1000",
   		34 => "0000",
   		35 => "0000",
   		36 => "1010",
   		37 => "1000",
   		38 => "0000",
   		39 => "0000",
   		40 => "1010",
   		41 => "1000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0010",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "1100",
   		50 => "0100",
   		51 => "0100",
   		52 => "1100",
   		53 => "1100",
   		54 => "0100",
   		55 => "0100",
   		56 => "1100",
   		57 => "1100",
   		58 => "0100",
   		59 => "0100",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0100",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 14
   constant routing_table_bits_14: t_tata_long := (
   	-- local
   		0 => "1000",
   		1 => "0000",
   		2 => "0000",
   		3 => "0000",
   		4 => "0000",
   		5 => "0000",
   		6 => "0000",
   		7 => "0000",
   		8 => "0000",
   		9 => "0000",
   		10 => "0000",
   		11 => "0000",
   		12 => "0000",
   		13 => "0000",
   		14 => "0000",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0000",
   		18 => "0000",
   		19 => "0000",
   		20 => "0000",
   		21 => "0000",
   		22 => "0000",
   		23 => "0000",
   		24 => "0000",
   		25 => "0000",
   		26 => "0000",
   		27 => "0000",
   		28 => "0000",
   		29 => "0000",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0010",
   		34 => "0000",
   		35 => "0000",
   		36 => "0010",
   		37 => "0010",
   		38 => "0000",
   		39 => "0000",
   		40 => "0010",
   		41 => "0010",
   		42 => "0000",
   		43 => "0000",
   		44 => "0010",
   		45 => "0010",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "0100",
   		50 => "0100",
   		51 => "0100",
   		52 => "0100",
   		53 => "0100",
   		54 => "0100",
   		55 => "0100",
   		56 => "0100",
   		57 => "0100",
   		58 => "0100",
   		59 => "0100",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0100",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );
   -- Node 15
   constant routing_table_bits_15: t_tata_long := (
   	-- local
   		0 => "0000",
   		1 => "1010",
   		2 => "1000",
   		3 => "1000",
   		4 => "1010",
   		5 => "1010",
   		6 => "1000",
   		7 => "1000",
   		8 => "1010",
   		9 => "1010",
   		10 => "1000",
   		11 => "1000",
   		12 => "0010",
   		13 => "0010",
   		14 => "0000",
   		15 => "0000",
   	-- north
   		16 => "0000",
   		17 => "0010",
   		18 => "0000",
   		19 => "0000",
   		20 => "0010",
   		21 => "0010",
   		22 => "0000",
   		23 => "0000",
   		24 => "0010",
   		25 => "0010",
   		26 => "0000",
   		27 => "0000",
   		28 => "0010",
   		29 => "0010",
   		30 => "0000",
   		31 => "0000",
   	-- east
   		32 => "0000",
   		33 => "0000",
   		34 => "0000",
   		35 => "0000",
   		36 => "0000",
   		37 => "0000",
   		38 => "0000",
   		39 => "0000",
   		40 => "0000",
   		41 => "0000",
   		42 => "0000",
   		43 => "0000",
   		44 => "0000",
   		45 => "0000",
   		46 => "0000",
   		47 => "0000",
   	-- west
   		48 => "0000",
   		49 => "1000",
   		50 => "1000",
   		51 => "1000",
   		52 => "1000",
   		53 => "1000",
   		54 => "1000",
   		55 => "1000",
   		56 => "1000",
   		57 => "1000",
   		58 => "1000",
   		59 => "1000",
   		60 => "0000",
   		61 => "0000",
   		62 => "0000",
   		63 => "0000",
   	-- south
   		64 => "0000",
   		65 => "0000",
   		66 => "0000",
   		67 => "0000",
   		68 => "0000",
   		69 => "0000",
   		70 => "0000",
   		71 => "0000",
   		72 => "0000",
   		73 => "0000",
   		74 => "0000",
   		75 => "0000",
   		76 => "0000",
   		77 => "0000",
   		78 => "0000",
   		79 => "0000"
    );



end type_def_pack;
